// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
// CREATED		"Fri Nov 26 14:42:59 2021"

module lab1(
	pin_name1,
	pin_name2,
	pin_name3,
	pin_name4,
	pin_name5,
	pin_name6,
	pin_name7,
	pin_name8,
	pin_name9,
	pin_name10,
	pin_name11,
	pin_name12,
	pin_name13,
	pin_name14,
	pin_name15,
	pin_name16,
	pin_name17,
	pin_name18,
	pin_name19,
	pin_name20,
	pin_name21,
	pin_name22,
	pin_name23,
	pin_name24
);


input wire	pin_name1;
input wire	pin_name2;
input wire	pin_name3;
input wire	pin_name4;
input wire	pin_name5;
input wire	pin_name6;
input wire	pin_name7;
input wire	pin_name8;
input wire	pin_name9;
input wire	pin_name10;
input wire	pin_name11;
input wire	pin_name12;
output wire	pin_name13;
output wire	pin_name14;
output wire	pin_name15;
output wire	pin_name16;
output wire	pin_name17;
output wire	pin_name18;
output wire	pin_name19;
output wire	pin_name20;
output wire	pin_name21;
output wire	pin_name22;
output wire	pin_name23;
output wire	pin_name24;


assign	pin_name13 = pin_name1;
assign	pin_name14 = pin_name2;
assign	pin_name15 = pin_name3;
assign	pin_name16 = pin_name4;
assign	pin_name17 = pin_name5;
assign	pin_name18 = pin_name6;
assign	pin_name19 = pin_name7;
assign	pin_name20 = pin_name8;
assign	pin_name21 = pin_name9;
assign	pin_name22 = pin_name10;
assign	pin_name23 = pin_name11;
assign	pin_name24 = pin_name12;




endmodule
